
module div_pll (
	refclk,
	rst,
	outclk_0,
	locked);	

	input		refclk;
	input		rst;
	output		outclk_0;
	output		locked;
endmodule
