
module pll50_25 (
	refclk,
	rst,
	outclk_0,
	locked);	

	input		refclk;
	input		rst;
	output		outclk_0;
	output		locked;
endmodule
