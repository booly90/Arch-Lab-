// div_pll.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module div_pll (
		output wire  locked,   //  locked.export
		output wire  outclk_0, // outclk0.clk
		input  wire  refclk,   //  refclk.clk
		input  wire  rst       //   reset.reset
	);

	div_pll_pll_0 pll_0 (
		.refclk   (refclk),   //  refclk.clk
		.rst      (rst),      //   reset.reset
		.outclk_0 (outclk_0), // outclk0.clk
		.locked   (locked)    //  locked.export
	);

endmodule
